module if (
    
);

endmodule 