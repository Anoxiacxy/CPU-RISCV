module stall_ctrl (
    input wire clk,
    input wire rst,

    input wire stall_if,
    input wire stall_id,
    input wire stall_ex,
    input wire stall_mem,

    output wire 
);
endmodule