module reg_id_ex (
    input wire clk,
    input wire rst,
    input wire [1 : 0] stall,

    

);
endmodule 