module icache (    
    input wire                  request,
    input wire [`MemAddrBus]    inst_addr,
    output reg                  inst_done,
    output reg [`MemDataBus]    inst_data,
);
endmodule